`timescale 1ns/1ps

module and_gate (
    input  logic a,
    input  logic b,
    output wire y   // <- cambiar a wire
);
    assign y = a & b;
endmodule
